library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
entity memory_rom is
	Port ( addr : in  STD_LOGIC_VECTOR (9 downto 0);
		output : out  STD_LOGIC_VECTOR (7 downto 0));
end memory_rom;

architecture Behavioral of memory_rom is
	type romtable is array (0 to 1023) of std_logic_vector(7 downto 0);

	constant romdata : romtable := (
		"00100110",
		"00010000",
		"01101111",
		"01110010",
		"00010010",
		"01111111",
		"01010111",
		"00000100",
		"00100101",
		"01000111",
		"01010100",
		"10010000",
		"11010001",
		"10110000",
		"01100110",
		"01100101",
		"10010101",
		"11010100",
		"01001101",
		"10111100",
		"10011001",
		"00001001",
		"00010001",
		"01000001",
		"00001011",
		"01100110",
		"11110100",
		"00000111",
		"11101011",
		"10111111",
		"00001111",
		"11100010",
		"10000001",
		"01100011",
		"11100000",
		"01000101",
		"11011001",
		"11100011",
		"00101101",
		"10111000",
		"10100010",
		"11011101",
		"10001010",
		"11101010",
		"00010110",
		"01100011",
		"01010101",
		"01111010",
		"11111011",
		"11111101",
		"00000010",
		"01011110",
		"10000111",
		"01010100",
		"11111001",
		"10111010",
		"11011011",
		"11110110",
		"00101110",
		"10111110",
		"00110011",
		"00001100",
		"00011111",
		"01010110",
		"10011101",
		"10100000",
		"00110000",
		"10110001",
		"00111100",
		"00000100",
		"11111011",
		"00000001",
		"01010110",
		"10011010",
		"10010101",
		"00101111",
		"00111010",
		"00110000",
		"00111101",
		"11001101",
		"11001000",
		"01101100",
		"11110100",
		"00010011",
		"11011011",
		"00010011",
		"00001100",
		"11111011",
		"01011111",
		"11111011",
		"11000000",
		"10110000",
		"10011100",
		"01010111",
		"01111011",
		"00001010",
		"01110010",
		"11110001",
		"10010100",
		"10000110",
		"00100000",
		"00100010",
		"01100100",
		"10010110",
		"00100100",
		"10100000",
		"01000001",
		"01000110",
		"10111101",
		"11111111",
		"01001010",
		"11000101",
		"11011000",
		"11010100",
		"10001100",
		"01000110",
		"01110101",
		"00001100",
		"10101111",
		"01110011",
		"10011011",
		"01100100",
		"11001111",
		"10010101",
		"11101010",
		"10001000",
		"00010101",
		"11010110",
		"00010011",
		"01100100",
		"01100110",
		"01110010",
		"01001100",
		"11011011",
		"10101000",
		"11100000",
		"10110111",
		"01011101",
		"11101101",
		"01101111",
		"00001111",
		"01110101",
		"11100011",
		"10110000",
		"00011111",
		"00001110",
		"00110000",
		"11110110",
		"11000110",
		"11000111",
		"10000001",
		"11010101",
		"00101000",
		"10001111",
		"11101110",
		"00001010",
		"00010111",
		"11111000",
		"11000010",
		"01011111",
		"10011100",
		"00110100",
		"00000100",
		"00011100",
		"10101010",
		"00100100",
		"01100111",
		"01010100",
		"11011111",
		"00000000",
		"11001111",
		"01010010",
		"01111011",
		"01101101",
		"11100011",
		"11000100",
		"01111001",
		"11011000",
		"11001110",
		"01000000",
		"10000000",
		"00110110",
		"01010110",
		"00100100",
		"10001001",
		"01010110",
		"01100000",
		"01011010",
		"11000010",
		"11110010",
		"10011011",
		"01010111",
		"10110010",
		"11111111",
		"11001001",
		"10010001",
		"01001100",
		"00101010",
		"11111101",
		"11011101",
		"00100000",
		"00010110",
		"10101111",
		"00011101",
		"10110000",
		"00100001",
		"11101111",
		"10101110",
		"11011011",
		"00101010",
		"11000001",
		"01110010",
		"11101110",
		"11001000",
		"11111101",
		"01001101",
		"10101100",
		"01111110",
		"00111101",
		"00010001",
		"00111001",
		"11000101",
		"01010110",
		"11111000",
		"00110101",
		"00111101",
		"00101001",
		"11001101",
		"10011000",
		"01100110",
		"10010001",
		"10011000",
		"01101100",
		"01000101",
		"00000000",
		"10100111",
		"00100100",
		"00101111",
		"00000001",
		"01001111",
		"10111101",
		"11110100",
		"10110110",
		"11100011",
		"11100100",
		"01100111",
		"00101010",
		"10010001",
		"11010010",
		"10100010",
		"00010101",
		"10000111",
		"01111011",
		"10110010",
		"11011010",
		"01010001",
		"11010101",
		"01001110",
		"01011101",
		"00010100",
		"00101111",
		"01010101",
		"00011001",
		"11010010",
		"00101011",
		"01100110",
		"10100011",
		"10110011",
		"10101001",
		"01100111",
		"10110011",
		"00010001",
		"01011001",
		"10011100",
		"11101010",
		"00110100",
		"00010011",
		"01010011",
		"11111110",
		"10111111",
		"01000100",
		"00001100",
		"01100001",
		"01010000",
		"11110101",
		"10101110",
		"10011011",
		"11111101",
		"01010001",
		"01001100",
		"10100001",
		"01010001",
		"11011010",
		"11000001",
		"00000010",
		"11010001",
		"10110010",
		"11011101",
		"10110001",
		"10110110",
		"00100001",
		"11000011",
		"10010011",
		"00111011",
		"00000011",
		"11111000",
		"01001110",
		"10100000",
		"00000110",
		"00100000",
		"10001100",
		"01101111",
		"11111011",
		"01101000",
		"00000100",
		"01000111",
		"11101010",
		"11001101",
		"11110010",
		"10001010",
		"10001000",
		"11100111",
		"01101010",
		"01001000",
		"01111100",
		"01000101",
		"01111000",
		"00010001",
		"11000001",
		"10100110",
		"00001001",
		"00010000",
		"10001110",
		"10010100",
		"00010000",
		"00111110",
		"01010110",
		"00101101",
		"11011000",
		"11101001",
		"11000100",
		"11011100",
		"01011010",
		"10000110",
		"01001010",
		"11100010",
		"11001110",
		"01100000",
		"00110010",
		"11001100",
		"00010100",
		"11011101",
		"11001000",
		"10000100",
		"10010011",
		"10001000",
		"10000011",
		"11110110",
		"01101110",
		"11100101",
		"11001110",
		"01110110",
		"00001100",
		"11010100",
		"00011100",
		"01110011",
		"00101100",
		"11110010",
		"01101101",
		"11011001",
		"01111000",
		"11111110",
		"00010011",
		"11001111",
		"01111110",
		"01100000",
		"00000111",
		"00101011",
		"10101000",
		"11011000",
		"00001011",
		"00110100",
		"11010111",
		"01101101",
		"10100010",
		"01100001",
		"11010110",
		"00011000",
		"11011101",
		"01001001",
		"10010100",
		"10001000",
		"00110110",
		"11101111",
		"10011001",
		"10100000",
		"01001110",
		"00011000",
		"01011000",
		"00000010",
		"01110010",
		"01111011",
		"11101111",
		"11010100",
		"01101001",
		"11011100",
		"11101000",
		"10011011",
		"10100110",
		"01100101",
		"11001001",
		"00010001",
		"01110010",
		"10001110",
		"01001111",
		"11001010",
		"11111001",
		"00111000",
		"00011111",
		"01100001",
		"11111101",
		"11011011",
		"11100010",
		"10011010",
		"10101110",
		"00100011",
		"10010100",
		"00111010",
		"01110001",
		"01110001",
		"10110110",
		"11101010",
		"10100111",
		"10010001",
		"11110010",
		"10010110",
		"10000111",
		"11011010",
		"00100000",
		"01110010",
		"01000111",
		"01010100",
		"11000100",
		"01101001",
		"10011101",
		"11110110",
		"01000010",
		"10101110",
		"01011010",
		"10101001",
		"10000101",
		"11101011",
		"01011111",
		"10100101",
		"10111000",
		"11101011",
		"10001111",
		"10111110",
		"10100110",
		"00000011",
		"00111101",
		"10011111",
		"01100001",
		"01101011",
		"01000111",
		"11001011",
		"11111000",
		"11000010",
		"11010101",
		"11001110",
		"00100001",
		"10110001",
		"00000101",
		"00111010",
		"00010000",
		"00110100",
		"01100110",
		"10100000",
		"00110011",
		"00000010",
		"10011110",
		"10010111",
		"11001111",
		"11111011",
		"01010011",
		"00011000",
		"10001110",
		"00001111",
		"11111010",
		"01111100",
		"10000100",
		"00010101",
		"11000100",
		"11000011",
		"01101011",
		"01001010",
		"00001100",
		"00110001",
		"10100010",
		"01110010",
		"01000001",
		"11011001",
		"00100110",
		"00100001",
		"00101110",
		"11100010",
		"01100010",
		"00101111",
		"00110111",
		"00100110",
		"00100000",
		"01011001",
		"00001111",
		"11000100",
		"11011010",
		"01111000",
		"00011000",
		"10011110",
		"01101001",
		"01011011",
		"00010101",
		"10011110",
		"01011011",
		"11110000",
		"01000011",
		"01000000",
		"10000101",
		"01001110",
		"01001011",
		"10100101",
		"10111110",
		"01000100",
		"00010010",
		"00000011",
		"10100000",
		"11000001",
		"11011111",
		"01100011",
		"00100010",
		"11010001",
		"11000010",
		"10010001",
		"00110011",
		"01001111",
		"01101111",
		"11001110",
		"10111001",
		"10101011",
		"11010101",
		"00101000",
		"11101110",
		"00010011",
		"11010000",
		"10000011",
		"10100000",
		"01101000",
		"10111100",
		"10001110",
		"01101100",
		"01010011",
		"10100101",
		"10100110",
		"00011010",
		"10110111",
		"10111110",
		"00101001",
		"00110011",
		"01110001",
		"00111011",
		"00100110",
		"10011111",
		"00000100",
		"11101001",
		"11111100",
		"10001100",
		"10011010",
		"10100101",
		"01110100",
		"10001000",
		"11101011",
		"00101101",
		"11110111",
		"10100001",
		"11001111",
		"11100111",
		"00101010",
		"01011000",
		"10001010",
		"11010011",
		"00100101",
		"01011011",
		"11101110",
		"01001110",
		"11010000",
		"10111000",
		"11010110",
		"11100001",
		"10111110",
		"00110110",
		"11111000",
		"01001101",
		"11000010",
		"00110011",
		"00010010",
		"11110100",
		"00000111",
		"00001111",
		"11010101",
		"01010010",
		"11011101",
		"00111000",
		"10011011",
		"11010111",
		"11001111",
		"10010011",
		"01111000",
		"11110001",
		"01110001",
		"00000000",
		"11111110",
		"01011001",
		"10010011",
		"01101101",
		"01011101",
		"00000110",
		"10110001",
		"00111000",
		"10100100",
		"10001000",
		"01000010",
		"01101000",
		"01101110",
		"11011011",
		"01000100",
		"01011000",
		"01010111",
		"10000000",
		"10011000",
		"00111111",
		"00001100",
		"10100100",
		"11101101",
		"00111000",
		"00001001",
		"11110111",
		"01000010",
		"00101101",
		"10111000",
		"11100111",
		"01100010",
		"10000011",
		"11001000",
		"11000010",
		"10110001",
		"00101100",
		"00011010",
		"10000101",
		"11101110",
		"11000000",
		"10100000",
		"01000000",
		"01010111",
		"00000001",
		"11110010",
		"11110110",
		"01101111",
		"11010011",
		"00000001",
		"11110010",
		"01010001",
		"10011101",
		"01101100",
		"11011101",
		"00000110",
		"10101011",
		"10000001",
		"10000000",
		"10111011",
		"01101110",
		"11011000",
		"11111110",
		"10011101",
		"01110110",
		"01100001",
		"11000110",
		"01110101",
		"00011011",
		"10110001",
		"10000100",
		"01100110",
		"10100001",
		"11111111",
		"01100100",
		"01000000",
		"00000011",
		"00110000",
		"11010010",
		"11011111",
		"10110110",
		"10010011",
		"01001110",
		"01000111",
		"11100001",
		"00101011",
		"01110000",
		"00001001",
		"11111101",
		"01110000",
		"11110110",
		"10010001",
		"11000010",
		"00100101",
		"11011010",
		"01100111",
		"01011111",
		"01100101",
		"10000100",
		"10011100",
		"00100010",
		"11000011",
		"10111000",
		"00110010",
		"00001000",
		"11011010",
		"00010000",
		"01001110",
		"01011110",
		"00010100",
		"10100100",
		"10100000",
		"11110010",
		"01100100",
		"10011000",
		"11111110",
		"00100101",
		"00111011",
		"01011000",
		"11100011",
		"00111000",
		"01111001",
		"11101111",
		"00101011",
		"11001001",
		"01011110",
		"00111001",
		"00110111",
		"01010000",
		"00111001",
		"01111101",
		"10101011",
		"11010010",
		"01101110",
		"00110011",
		"00110101",
		"00100000",
		"10011010",
		"00100000",
		"01100101",
		"11111001",
		"00010111",
		"11101100",
		"10011001",
		"10010000",
		"10111100",
		"00011110",
		"10000010",
		"00100101",
		"10101101",
		"11010011",
		"01100100",
		"11110111",
		"10101011",
		"10010100",
		"11010111",
		"00110001",
		"00010101",
		"10010011",
		"10001111",
		"00000110",
		"11011000",
		"10010101",
		"10101101",
		"10101100",
		"00111100",
		"10111111",
		"10101101",
		"01110101",
		"01011010",
		"00001110",
		"10010000",
		"01100110",
		"10100001",
		"00111011",
		"00000000",
		"10111000",
		"01010100",
		"11011101",
		"10000001",
		"01000000",
		"01100101",
		"00010011",
		"01101010",
		"10010000",
		"11011111",
		"11110010",
		"10100000",
		"00111110",
		"10001110",
		"00000111",
		"10000001",
		"11001100",
		"10001110",
		"01000101",
		"10100111",
		"11100000",
		"00001101",
		"00000001",
		"01101000",
		"11001000",
		"00010010",
		"01101101",
		"01110111",
		"11101101",
		"00100001",
		"11100111",
		"10010001",
		"10111001",
		"01111000",
		"11001110",
		"01101111",
		"10010001",
		"00010001",
		"10100000",
		"01011100",
		"10101011",
		"01001010",
		"11111111",
		"11100101",
		"00110000",
		"10001110",
		"00101010",
		"10010100",
		"10110110",
		"11000101",
		"11111010",
		"10111010",
		"00101000",
		"11110100",
		"11100011",
		"00010110",
		"10100101",
		"01111110",
		"10010101",
		"00001010",
		"00011000",
		"01111010",
		"01101111",
		"10100000",
		"00100000",
		"11101001",
		"01110101",
		"11110110",
		"11001000",
		"10100110",
		"11110111",
		"10010111",
		"00110000",
		"01000011",
		"10110001",
		"00001100",
		"11101101",
		"00010101",
		"11011000",
		"00000001",
		"01111111",
		"01000101",
		"00101101",
		"00101111",
		"11000110",
		"00101101",
		"11100100",
		"01011000",
		"10010100",
		"11100101",
		"01001011",
		"11001000",
		"00000011",
		"10011001",
		"10100010",
		"01011100",
		"10010111",
		"11001010",
		"11111011",
		"00111110",
		"10011101",
		"00110111",
		"00111011",
		"00011000",
		"00111101",
		"10011111",
		"00010101",
		"10000000",
		"01010001",
		"00110000",
		"01100110",
		"10000101",
		"00011101",
		"11111111",
		"00011111",
		"11100111",
		"01010000",
		"01111111",
		"11010100",
		"11010100",
		"00111011",
		"10001101",
		"00010011",
		"11010100",
		"11101011",
		"10101110",
		"01101010",
		"11010010",
		"11011000",
		"01111011",
		"00110001",
		"10000001",
		"10000010",
		"00010100",
		"01001000",
		"00000011",
		"10010100",
		"10111101",
		"00010000",
		"00011100",
		"10101100",
		"10011000",
		"00100101",
		"00011011",
		"10100111",
		"11011111",
		"10100110",
		"11101010",
		"00100001",
		"10001111",
		"00101000",
		"11001011",
		"00000001",
		"00100010",
		"00010011",
		"11101010",
		"01001010",
		"10010110",
		"11111000",
		"01010110",
		"10100001",
		"10011100",
		"01110110",
		"11111110",
		"10011110",
		"11111111",
		"11110011",
		"00011010",
		"01010110",
		"01110011",
		"10000110",
		"00110000",
		"00001101",
		"01110001",
		"01100110",
		"10011011",
		"01111001",
		"11011111",
		"00001110",
		"11101111",
		"01011010",
		"01010110",
		"11110011",
		"11000110",
		"01011101",
		"00111010",
		"10110101",
		"00100000",
		"10011000",
		"01111010",
		"11110010",
		"00001010",
		"11101001",
		"11010111",
		"01001101",
		"00011110",
		"01011100",
		"00101110",
		"00011101",
		"10001001",
		"11000000",
		"00101001",
		"00001011",
		"10100001",
		"10111111",
		"10101111",
		"01110101",
		"10110101",
		"01010100",
		"00011001",
		"10111100",
		"10111101",
		"00000100",
		"11101100",
		"11000000",
		"01100010",
		"00101100",
		"01011000",
		"10100101",
		"11111000",
		"01010111",
		"00010000",
		"01010001",
		"11111110",
		"01100111",
		"10010011",
		"11001011",
		"10001101",
		"00011100",
		"10101110"
		);

begin
  process (addr)
  begin
		output <= romdata (conv_integer(addr));
  end process;
end Behavioral;
